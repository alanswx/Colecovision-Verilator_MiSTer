
module cv_adamnet (
  input        clk_i,
  input        adam_reset_pcb_n_i /*verilator public_flat*/,
  input        z80_wr/*verilator public_flat*/,
  input        z80_rd/*verilator public_flat*/,
  input [15:0] z80_addr/*verilator public_flat*/,
  input [7:0]  z80_data/*verilator public_flat*/
);



endmodule
